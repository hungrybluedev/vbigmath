module main

import big
import crypto.sha1
import rand

fn main() {
	// zm := _000
	zs := 20_000

	rand.seed([u32(314981), 1397])

	for _ in 0 .. 20 {
		x, y := zs, zs
		z := x + y

		a1, a2 := rand.int_in_range(1, 101)?, rand.int_in_range(1, 101)?

		b1 := big.integer_from_string(a1.str() + '0'.repeat(x))?
		b2 := big.integer_from_string(a2.str() + '0'.repeat(y))?

		c := b1 * b2
		c_str := c.str()
		assert c_str == (a1 * a2).str() + '0'.repeat(z)
		println(sha1.hexhash(c_str) + ' ' + (c.bit_len() / 32).str())
	}
	// values := [
	// 	// [
	// 	// 	'4198374698153841387469138475139192391476981638148746183691874647987364918736498713694879861387463981734698173469813746918734613987416898173498369131982649871694871364133413987469238476193874691837469183746918374698137469813746981345987134689137569831746998371569837650398476982734693847058692874631987461938491873141',
	// 	// 	'1049861087364918641625457851369817346987136491387548715188691834419874698165936459419238716951498370197569138478013984769183649137468917349693769183746187416387469816350958734659832750937865098345709348537245609384560392744444444295602348307945603478509832709657160975098345607651301091650371614861938745193654913414',
	// 	// ],
	// 	[
	// 		'18746138746987365987519872364189480172146019374691864501346103786491387560138465103847017354360401387460183745183746103874613603178516036503465138746031874658361501378460139746836017346071356081371074613974603501387461374601378461350137461039746013974601738560137460173409138746013746873156137460134710378461387610344',
	// 		'1049861087364918641625457851369817346987136491387548715188691834419874698165936459419238716951498370197569138478013984769183649137468917349693769183746187416387469816350958734659832750937865098345709348537245609384560392744444444295602348307945603478509832709657160975098345607651301091650371614861938745193654913414',
	// 	],
	// 	// ['123', '456']
	// ]

	// for p in values {
	// 	a := big.integer_from_string(p[0])?
	// 	b := big.integer_from_string(p[1])?

	// 	println(a * b)
	// }
}
